module IR_FSM_bak(
			sysclk,
			reset,
			IRData,
			
			SegData,
			StoreCode,
			FushCode

);

input wire sysclk;
input wire reset;
input wire[31:0] IRData;

output wire[31:0] SegData;
output wire 		StoreCode;
output wire 		FushCode;







endmodule