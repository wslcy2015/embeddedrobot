module SW(
			sw,
			seg,
			binary
);

input [17:0] sw;

output reg [11:0] seg;
output reg [8:0] 	binary;

